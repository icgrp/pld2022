module bft_level_0(
  input clk,
  input [195:0] din0,
  input [195:0] din1,
  input [195:0] din2,
  input [195:0] din3,
  input reset,
  output [195:0] l_bus_o,
  output [195:0] l_but_o1,
  output [195:0] r_but_o,
  output [195:0] r_but_o1);



endmodule
