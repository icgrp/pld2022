module bft(
  input clk,
  input reset,
  input [48:0]dout_leaf_0,
  input [48:0]dout_leaf_1,
  input [48:0]dout_leaf_2,
  input [48:0]dout_leaf_3,
  input [48:0]dout_leaf_4,
  input [48:0]dout_leaf_5,
  input [48:0]dout_leaf_6,
  input [48:0]dout_leaf_7,
  input [48:0]dout_leaf_8,
  input [48:0]dout_leaf_9,
  input [48:0]dout_leaf_10,
  input [48:0]dout_leaf_11,
  input [48:0]dout_leaf_12,
  input [48:0]dout_leaf_13,
  input [48:0]dout_leaf_14,
  input [48:0]dout_leaf_15,
  input [48:0]dout_leaf_16,
  input [48:0]dout_leaf_17,
  input [48:0]dout_leaf_18,
  input [48:0]dout_leaf_19,
  input [48:0]dout_leaf_20,
  input [48:0]dout_leaf_21,
  input [48:0]dout_leaf_22,
  input [48:0]dout_leaf_23,
  input [48:0]dout_leaf_24,
  input [48:0]dout_leaf_25,
  input [48:0]dout_leaf_26,
  input [48:0]dout_leaf_27,
  input [48:0]dout_leaf_28,
  input [48:0]dout_leaf_29,
  input [48:0]dout_leaf_30,
  input [48:0]dout_leaf_31,
  output [48:0]din_leaf_0,
  output [48:0]din_leaf_1,
  output [48:0]din_leaf_2,
  output [48:0]din_leaf_3,
  output [48:0]din_leaf_4,
  output [48:0]din_leaf_5,
  output [48:0]din_leaf_6,
  output [48:0]din_leaf_7,
  output [48:0]din_leaf_8,
  output [48:0]din_leaf_9,
  output [48:0]din_leaf_10,
  output [48:0]din_leaf_11,
  output [48:0]din_leaf_12,
  output [48:0]din_leaf_13,
  output [48:0]din_leaf_14,
  output [48:0]din_leaf_15,
  output [48:0]din_leaf_16,
  output [48:0]din_leaf_17,
  output [48:0]din_leaf_18,
  output [48:0]din_leaf_19,
  output [48:0]din_leaf_20,
  output [48:0]din_leaf_21,
  output [48:0]din_leaf_22,
  output [48:0]din_leaf_23,
  output [48:0]din_leaf_24,
  output [48:0]din_leaf_25,
  output [48:0]din_leaf_26,
  output [48:0]din_leaf_27,
  output [48:0]din_leaf_28,
  output [48:0]din_leaf_29,
  output [48:0]din_leaf_30,
  output [48:0]din_leaf_31,
  output resend_0,
  output resend_1,
  output resend_2,
  output resend_3,
  output resend_4,
  output resend_5,
  output resend_6,
  output resend_7,
  output resend_8,
  output resend_9,
  output resend_10,
  output resend_11,
  output resend_12,
  output resend_13,
  output resend_14,
  output resend_15,
  output resend_16,
  output resend_17,
  output resend_18,
  output resend_19,
  output resend_20,
  output resend_21,
  output resend_22,
  output resend_23,
  output resend_24,
  output resend_25,
  output resend_26,
  output resend_27,
  output resend_28,
  output resend_29,
  output resend_30,
  output resend_31);
    // empty
    gen_nw32 # (
        .num_leaves(32),
        .payload_sz(43),
        .p_sz(49),
        .addr(1'b0),
        .level(0)
        ) gen_nw32 (
        .clk(clk),
        .reset(reset),
        .pe_interface(
            {
            dout_leaf_31,
            dout_leaf_30,
            dout_leaf_29,
            dout_leaf_28,
            dout_leaf_27,
            dout_leaf_26,
            dout_leaf_25,
            dout_leaf_24,
            dout_leaf_23,
            dout_leaf_22,
            dout_leaf_21,
            dout_leaf_20,
            dout_leaf_19,
            dout_leaf_18,
            dout_leaf_17,
            dout_leaf_16,
            dout_leaf_15,
            dout_leaf_14,
            dout_leaf_13,
            dout_leaf_12,
            dout_leaf_11,
            dout_leaf_10,
            dout_leaf_9,
            dout_leaf_8,
            dout_leaf_7,
            dout_leaf_6,
            dout_leaf_5,
            dout_leaf_4,
            dout_leaf_3,
            dout_leaf_2,
            dout_leaf_1,
            dout_leaf_0}),
        .interface_pe(
            {
           din_leaf_31,
           din_leaf_30,
           din_leaf_29,
           din_leaf_28,
           din_leaf_27,
           din_leaf_26,
           din_leaf_25,
           din_leaf_24,
           din_leaf_23,
           din_leaf_22,
           din_leaf_21,
           din_leaf_20,
           din_leaf_19,
           din_leaf_18,
           din_leaf_17,
           din_leaf_16,
           din_leaf_15,
           din_leaf_14,
           din_leaf_13,
           din_leaf_12,
           din_leaf_11,
           din_leaf_10,
           din_leaf_9,
           din_leaf_8,
           din_leaf_7,
           din_leaf_6,
           din_leaf_5,
           din_leaf_4,
           din_leaf_3,
           din_leaf_2,
           din_leaf_1,
           din_leaf_0}),
        .resend(
            {
            resend_31,
            resend_30,
            resend_29,
            resend_28,
            resend_27,
            resend_26,
            resend_25,
            resend_24,
            resend_23,
            resend_22,
            resend_21,
            resend_20,
            resend_19,
            resend_18,
            resend_17,
            resend_16,
            resend_15,
            resend_14,
            resend_13,
            resend_12,
            resend_11,
            resend_10,
            resend_9,
            resend_8,
            resend_7,
            resend_6,
            resend_5,
            resend_4,
            resend_3,
            resend_2,
            resend_1,
            resend_0})
    );
endmodule
